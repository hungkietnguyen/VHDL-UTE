----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:27:31 04/08/2023 
-- Design Name: 
-- Module Name:    LCD_GAN_DULIEU_GPG_NN - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity LCD_GAN_DULIEU_GPG_NN is
    Port ( GT_MOD : in  STD_LOGIC_VECTOR (1 downto 0);
           DV_GIAY : in  STD_LOGIC_VECTOR (3 downto 0);
           CH_GIAY : in  STD_LOGIC_VECTOR (3 downto 0);
           DV_PHUT : in  STD_LOGIC_VECTOR (3 downto 0);
           CH_PHUT : in  STD_LOGIC_VECTOR (3 downto 0);
           DV_GIO : in  STD_LOGIC_VECTOR (3 downto 0);
           CH_GIO : in  STD_LOGIC_VECTOR (3 downto 0);
           
			  ENA2HZ : in  STD_LOGIC;
           CD_BUP : in  STD_LOGIC;
           CD_BDW : in  STD_LOGIC;
           CKHT : in  STD_LOGIC;
			  ND_TR : in  STD_LOGIC_VECTOR (3 downto 0);
			  ND_CH : in  STD_LOGIC_VECTOR (3 downto 0);
			  ND_DV : in  STD_LOGIC_VECTOR (3 downto 0);
           DA_TR : in  STD_LOGIC_VECTOR (3 downto 0);
			  DA_CH : in  STD_LOGIC_VECTOR (3 downto 0);
			  DA_DV : in  STD_LOGIC_VECTOR (3 downto 0);
			  TT_CS,DHT_PR:  in  STD_LOGIC;
           LCD_H0 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_H1 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_H2 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_H3 : out  STD_LOGIC_VECTOR (159 downto 0));
end LCD_GAN_DULIEU_GPG_NN;

architecture Behavioral of LCD_GAN_DULIEU_GPG_NN is
SIGNAL DVGIO_NN : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DVPHUT_NN : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DVGIAY_NN : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL CHGIO_NN : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL CHPHUT_NN : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL CHGIAY_NN : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL Q_R, Q_N :STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL DHT0,DHT1,DHT2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
begin
	PROCESS(DHT_PR,TT_CS)
	BEGIN 
		IF (DHT_PR='1') THEN
			DHT2<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
			DHT1<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
			DHT0<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
		ELSIF(TT_CS='0') THEN
			DHT2<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
			DHT1<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
			DHT0<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8);
		ELSE	
			DHT2<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
			DHT1<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
			DHT0<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
		END IF;
	END PROCESS;
	
	PROCESS(CKHT)
	BEGIN 
		IF FALLING_EDGE(CKHT) THEN Q_R <= Q_N;
		END IF;
	END PROCESS;
	
	PROCESS(CKHT)
	BEGIN 
		IF FALLING_EDGE(CKHT) THEN Q_R <= Q_N;
		END IF;
	END PROCESS;
	
	PROCESS(Q_R,GT_MOD,ENA2HZ,CD_BUP,CD_BDW)
	BEGIN
		Q_N <= Q_R;
		 IF ENA2HZ ='1' THEN
			IF CD_BUP ='0' AND CD_BDW ='0' THEN
				IF GT_MOD ="01" THEN Q_N <="11" & NOT Q_R(0);
				ELSIF GT_MOD="10" THEN Q_N <= '1' & NOT Q_R(1) &'1';
				ELSIF GT_MOD="11" THEN Q_N <= NOT Q_R(2) & "11";
				ELSE  Q_N <= "111" ;
				END IF;
			ELSE Q_N <= "111";	
			END IF;
		END IF;
	END PROCESS;
	CHGIO_NN <= X"3" & CH_GIO WHEN Q_R(2) ='1' ELSE X"20";
	DVGIO_NN <= X"3" & DV_GIO WHEN Q_R(2) ='1' ELSE X"20";
	
	CHPHUT_NN <= X"3" & CH_PHUT WHEN Q_R(1) ='1' ELSE X"20";
	DVPHUT_NN <= X"3" & DV_PHUT WHEN Q_R(1) ='1' ELSE X"20";
	
	CHGIAY_NN <= X"3" & CH_GIAY WHEN Q_R(0) ='1' ELSE X"20";
	DVGIAY_NN <= X"3" & DV_GIAY WHEN Q_R(0) ='1' ELSE X"20";
--HANG 0	
	 LCD_H0( 7 DOWNTO 0)     <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	 LCD_H0(15 DOWNTO 8)   	 <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('L'),8);
	 LCD_H0(23 DOWNTO 16)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	 LCD_H0(31 DOWNTO 24)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	 LCD_H0(39 DOWNTO 32)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	 LCD_H0(47 DOWNTO 40)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	 LCD_H0(55 DOWNTO 48)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('G'),8);
	 LCD_H0(63 DOWNTO 56)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('P'),8);
	 LCD_H0(71 DOWNTO 64)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('G'),8);
	 LCD_H0(79 DOWNTO 72)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	 LCD_H0(87 DOWNTO 80)    <= X"3" & "00"& GT_MOD;
	 LCD_H0(95 DOWNTO 88)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	 
	 LCD_H0(103 DOWNTO 96)   <= CHGIO_NN;
	 LCD_H0(111 DOWNTO 104)  <= DVGIO_NN;
	 LCD_H0(119 DOWNTO 112)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('-'),8);
	 LCD_H0(127 DOWNTO 120)  <= CHPHUT_NN;
	 LCD_H0(135 DOWNTO 128)  <= DVPHUT_NN;
	
	 LCD_H0(143 DOWNTO 136) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('-'),8);
	 LCD_H0(151 DOWNTO 144) <= CHGIAY_NN;
	 LCD_H0(159 DOWNTO 152) <= DVGIAY_NN;
---HANG 1	 
	 LCD_H1(7 DOWNTO 0)      <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
	 LCD_H1(15 DOWNTO 8)   	 <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	 LCD_H1(23 DOWNTO 16)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	 LCD_H1(31 DOWNTO 24)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	 LCD_H1(39 DOWNTO 32)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	 LCD_H1(47 DOWNTO 40)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	 LCD_H1(55 DOWNTO 48)    <= DHT2;
	 LCD_H1(63 DOWNTO 56)    <= DHT1;
	 LCD_H1(71 DOWNTO 64)    <= DHT0;
	 LCD_H1(79 DOWNTO 72)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	 LCD_H1(87 DOWNTO 80)    <= X"20" WHEN ND_TR=X"0" ELSE X"3" &ND_TR;
	 LCD_H1(95 DOWNTO 88)    <= X"3" &ND_CH;
	 LCD_H1(103 DOWNTO 96)   <= X"3" &ND_DV;
	 LCD_H1(111 DOWNTO 104)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	 LCD_H1(119 DOWNTO 112)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
	 LCD_H1(127 DOWNTO 120)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	 LCD_H1(135 DOWNTO 128)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	 LCD_H1(143 DOWNTO 136)  <= X"20" WHEN DA_TR=X"0" ELSE X"3" &DA_TR;
	 LCD_H1(151 DOWNTO 144)  <= X"3" &DA_CH;
	 LCD_H1(159 DOWNTO 152)  <= X"3" &DA_DV;
--HANG2	 
	 LCD_H2(7 DOWNTO 0)      <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	 LCD_H2(15 DOWNTO 8)   	 <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	 LCD_H2(23 DOWNTO 16)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('I'),8);
	 LCD_H2(31 DOWNTO 24)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8);
	 LCD_H2(39 DOWNTO 32)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	 LCD_H2(47 DOWNTO 40)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	 LCD_H2(55 DOWNTO 48)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	 LCD_H2(63 DOWNTO 56)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8);
	 LCD_H2(71 DOWNTO 64)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	 LCD_H2(79 DOWNTO 72)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('V'),8);
	 LCD_H2(87 DOWNTO 80)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('I'),8);
	 LCD_H2(95 DOWNTO 88)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	 LCD_H2(103 DOWNTO 96)   <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('M'),8);
	 LCD_H2(111 DOWNTO 104)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	 LCD_H2(119 DOWNTO 112)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	 LCD_H2(127 DOWNTO 120)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	 LCD_H2(135 DOWNTO 128)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	 LCD_H2(143 DOWNTO 136)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('S'),8);
	 LCD_H2(151 DOWNTO 144)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	 LCD_H2(159 DOWNTO 152)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
--HANG3	 
	 LCD_H3(7 DOWNTO 0)      <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
	 LCD_H3(15 DOWNTO 8)   	 <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	 LCD_H3(23 DOWNTO 16)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('I'),8);
	 LCD_H3(31 DOWNTO 24)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	 LCD_H3(39 DOWNTO 32)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	 LCD_H3(47 DOWNTO 40)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('F'),8);
	 LCD_H3(55 DOWNTO 48)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('P'),8);
	 LCD_H3(63 DOWNTO 56)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('G'),8);
	 LCD_H3(71 DOWNTO 64)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	 LCD_H3(79 DOWNTO 72)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	 LCD_H3(87 DOWNTO 80)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('X'),8);
	 LCD_H3(95 DOWNTO 88)    <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	 LCD_H3(103 DOWNTO 96)   <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('3'),8);
	 LCD_H3(111 DOWNTO 104)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('S'),8);
	 LCD_H3(119 DOWNTO 112)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('5'),8);
	 LCD_H3(127 DOWNTO 120)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('0'),8);
	 LCD_H3(135 DOWNTO 128)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('0'),8);
	 LCD_H3(143 DOWNTO 136)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8);
	 LCD_H3(151 DOWNTO 144)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
	 LCD_H3(159 DOWNTO 152)  <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
 
end Behavioral;

